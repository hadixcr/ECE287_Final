//module to detect when sound occurs in an audio file. 
module sound_analyzer();